DMM_AC_TO_DC1.CIR
*
* INPUT VOLTAGE
VIN	1	0	SIN(0V 1V 60HZ)
*
* RC INPUT
C1	1	2	10UF
R1	2	3	10k
*
* AMP AND DC FEEDBACK
XOP1	0 3 4	OPAMP1
RDC1	3	7	10K
CDC1	7	0	10UF
RDC2	7	4	10K
* POS CYCLE
R2		3	5	10K
R3		5	0	2K
D1		4	5	D1N4148
*
*  NEG CYCLE
R4		3	6	10K
R5		6	0	2K
D2		6	4	D1N4148
*
* LOW PASS FILTER
RLP1	5	8	100K
CLP1	0	0	1UF
RLP2	8	9	100K
CLP2	9	0	1UF

*
* DIODE
.model	D1N4148	D(Is=0.1p Rs=16 CJO=2p Tt=12n Bv=100 Ibv=0.1p)
*
* OPAMP MACRO MODEL, SINGLE-POLE *********
*
* connections:      +   -   out
.SUBCKT OPAMP1	    1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
EGAIN	3 0	1 2	100K
RP1	3	4	100K
CP1	4	0	0.159UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS
*
* ANALYSIS *************************************************
*.TRAN 	10US  100MS
.TRAN 	10US  1000MS 900MS

.control
run
plot v(1) v(9)
.endc

.END
