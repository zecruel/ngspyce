* teste da geracao de CM -> filtro media movel

* .---------------------------------.
* | Descricao do circuito principal |
* `---------------------------------'
vent 2 1 dc 0 sin(0 1 1k)
vruido 1 0 dc 0 trnoise(0.2 1e-5 0 0) ;ruido branco, ampl = 0.2, amostr = 10us
afilt 2 3 filtro
rzin 2 0 10k
rsaida 3 0 10k

* .--------------------------.
* | Descricao de componentes |
* `--------------------------'
.model filtro sma(pontos = 20, passo = 1e-5)

* .--------------------------------------.
* | Parametros de analise de Transitorio |
* `--------------------------------------'
*ATENCAO: Sempre considerar as condicoes iniciais (parametro uic)
*passo de amostragem = 10us, tempo total de 4ms
.tran 1e-5 4e-3 uic

* .------------------------------------.
* | Bloco de controle do Interpretador |
* `------------------------------------'
.control
run ; executa a simulacao
plot v(3) v(2)

*wrdata teste.txt v(node1) ; salva o resultado da simulacao em teste.txt
*quit ;sai do programa
.endc

* .--------------------------------------.
* |             ---- FIM ---             |
* `--------------------------------------'
.end