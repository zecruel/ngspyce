OP_PID1.CIR - OPAMP PID CONTROLLER
*
* SET POINT
VSET	1	0	PWL(0MS 0MV   0.1MS 0.1V   2000MS 0.1V)
*
* CALCULATE ERROR
R1	1	3	10K
R2	0	3	10K
R3	3	4	10K
XOP1	0 3 4	OPAMP1
*
* P - PROPORTIONAL TERM
RP1	4	5	1K
RP2	5	6	2K
XOP2	0 5 6	OPAMP1
*
* D - DERIVATIVE TERM
CD	4	7	0.1UF
RC	7	8	200
RD	8	9	1K
XOP3	0 8 9	OPAMP1
*
* I - INTEGRAL TERM
RI	4	10	100MEG
CI	10	11	1UF IC=0
XOP4	0 10 11	OPAMP1
*
* SIM PID TERMS
R4	6	12	10K
R5	9	12	10K
R6	11	12	10K
R7	12	13	10K
XOP5	0 12 13	OPAMP1
*
* INVERT SUMMATION
R8	13	14	10K
R9	14	15	10K
XOP6	0 14 15	OPAMP1
*
* PROCESS BLOCK WITH TIME LAG (PHASE SHIFT)
EOUT	20 0	15 0	100
RL1	20	21	10K
CL1	21	0	1UF
RL2	21	22	10K
CL2	22	0	1UF
*
* SENSOR BLOCK (NEG OUT FOR ERROR AMP.)
ESENSOR	23 0	22 0	-0.01
RL3	23	0	10K
*
* OPAMP MACRO MODEL, SINGLE-POLE WITH 10V OUTPUT CLAMP
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1	    1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN=100K AND POLE1=100HZ
* UNITY GAIN = DCGAIN X POLE1 = 10MHZ
EGAIN	3 0	1 2	100K
RP1	3	4	100K
CP1	4	0	0.0159UF
* ZENER LIMITER 
D1	4	7	DZ
D2	0	7	DZ
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
*
.model	DZ	D(Is=0.05u Rs=0.1 Bv=10 Ibv=0.05u)
.ENDS
*
* ANALYSIS
.TRAN 	0.1MS 10MS
*
* VIEW RESULTS
.PRINT TRAN	V(23)
.PROBE
.END