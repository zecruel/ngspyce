* teste da geracao de CM
vin 1 0 sin(0 1 1k)
ccouple 1 in 10uF
rzin in 0 19.35k

aamp in aout gain_block

rzout aout coll 3.9k
rbig coll 0 1e12

.model gain_block ganho(gain = -3.9 out_offset = 7.003)
.tran 1e-5 2e-3
.end